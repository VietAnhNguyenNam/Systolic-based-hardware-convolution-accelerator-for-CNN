--library IEEE;
--use IEEE.STD_LOGIC_1164.ALL;
--use IEEE.NUMERIC_STD.ALL;
--use work.common.all;

--entity Core is
--  generic (
--    B             : integer      := hyperparam_B;
--    K             : integer      := hyperparam_K;
--    BIAS_WIDTH    : integer      := hyperparam_BIAS_WIDTH;
--    MUX_SIZE      : integer      := hyperparam_MUX_SIZE;
--    MUX_SEL_WIDTH : integer      := hyperparam_MUX_SEL_WIDTH;
--    SB_LEN        : SB_len_t     := hyperparam_SB_LEN;
--    LEAFNO        : integer      := hyperparam_K;
--    LEAF_WIDTH    : integer      := hyperparam_LEAF_WIDTH;
--    ROOT_WIDTH    : integer      := hyperparam_SLICE_TREE_ROOT_WIDTH;
    
--    P_M           : integer      := hyperparam_P_M
--  );
--  port (
----    I_ext : in 
--  );
--end Core;

--architecture rtl of Core is

--begin


--end rtl;
